library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- decoder used in the registre file

entity decoder3_8 is
	port(
		regSlt : in std_logic_vector(4 downto 0);
		regOut : out std_logic
	);
	
end entity decoder3_8;

architecture RTL of decoder3_8 is
	
begin

end architecture RTL;
