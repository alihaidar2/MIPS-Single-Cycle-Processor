--Architecture------------	
begin
	
		outerloop: for i in 0 to 31 generate

--Most significant bit of aluOP (aluOP(2)) will determine Cin for add/sub operation. Cin=1 for sub
-- Set the initial Cin to 1 instead of 0, thus adding an extra 1 to the sum	for a sub operation	
		innerloop1: if (i = 0) generate
			addSub0: add_sub port map(Cin => aluOP(2), x => aluIn1(i), y => aluIn2(i),
										s => sig_aluOut(i), Cout => carry(i));
		end generate innerloop1;
		
		innerloop2: if (i>0 and i<31) generate 
				addsub: add_sub port map(Cin => carry(i-1), x => aluIn1(i), y => aluIn2(i),
										s => sig_aluOut(i), Cout => carry(i));
		end generate innerloop2;
		
		innerloop3: if (i=31) generate
			add31: add_sub port map (Cin => carry(i-1), x => aluIn1(i), y => aluIn2(i),
										s => sig_aluOut(i), Cout => CarryOut);
		end generate innerloop3;
		
	end generate outerloop;
	
	overflow: ofDetector port map(a => aluIn1(31), b => aluIn2(31), result => sig_aluOut(31), ovrflw => ovrflw);
	operation: mux32x4 port map(sel => aluOP(1 downto 0), logicAND => sig_AND, logicOR => sig_OR, add_sub => sig_aluOut, 
									SLT => sig_SLT, z => aluOut);

	sig_OR <= aluIn1 or aluIn2;
	sig_AND <= aluIn1 and aluIn2;
	
	zero <= not(sig_aluOut(0) or sig_aluOut(1) or sig_aluOut(2) or sig_aluOut(3) or sig_aluOut(4) or sig_aluOut(5) or
		 sig_aluOut(6) or sig_aluOut(7) or sig_aluOut(8) or sig_aluOut(9) or sig_aluOut(10) or sig_aluOut(11) or sig_aluOut(12) or
		  sig_aluOut(13) or sig_aluOut(14) or sig_aluOut(15) or sig_aluOut(16) or sig_aluOut(17) or sig_aluOut(18) or sig_aluOut(19) or
		   sig_aluOut(20) or sig_aluOut(21) or sig_aluOut(22) or sig_aluOut(23) or sig_aluOut(24) or sig_aluOut(25) or sig_aluOut(26) or
		    sig_aluOut(27) or sig_aluOut(28) or sig_aluOut(29) or sig_aluOut(30) or sig_aluOut(31));
		    	
	sig_SLT(31 downto 1) <= (others=>'0');
	sig_SLT(0) <= sig_aluOut(31); --For the least significant bit, SLT value should be sign of (aluIn1 - aluIn2)
	
end architecture;	

-- Linking of components and top level entity-----------
configuration conf_aluMain of aluMain is
	for aluMainArch
		for all : add_sub
			use entity work.add_sub(behave);
		end for;
		for all : ofDetector
			use entity work.ofDetector(behave);
		end for;
		for all : mux32x4
			use entity work.mux32x4(muxBehave);
		end for;
	end for;
end conf_aluMain;	
	
	
	
